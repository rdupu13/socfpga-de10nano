library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mantissa_unit is
	port
	(
		clk : in std_logic;
		rst : in std_logic
	);
end entity;

architecture mantissa_arch of mantissa is
	
	
	
	begin
		
		
		
end architecture;
