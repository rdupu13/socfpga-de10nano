library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity exponent_unit is
	port
	(
		clk : in  std_logic;
		rst : in  std_logic;
	
	);
end entity;

architecture exponent_unit_arch of exponent_unit is
	
	
	
	begin
		
		
		
end architecture;
